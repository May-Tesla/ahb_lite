
`ifndef AHB_DEFINE
    `define AHB_DEFINE

    `define IDLE   2'b00
    `define BUSY   2'b01
    `define NONSEQ 2'b10
    `define SEQ    2'b11
    
    `define SINGLE 3'b000
    `define INCR   3'b001
    `define WRAP4  3'b010
    `define INCR4  3'b011
    `define WRAP8  3'b100
    `define INCR8  3'b101
    `define WRAP16 3'b110
    `define INCR16 3'b111
    
    `define OKAY  2'b00
    `define ERROR 2'b01

`endif